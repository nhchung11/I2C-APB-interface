module i2c_core
(
	input wire          clk,
	input wire          rst_n,
    input wire          enable,
	input wire [6:0]    slave_address,
    input wire [7:0]    data_in,
    input wire          rw,
    input               sda_i, scl_i,
    output              sda_o, scl_o
	// inout               sda,        // tristate
	// inout               scl         // tristate
);

// FSM
localparam IDLE =           3'b000;
localparam START =          3'b001;
localparam WRITE_ADDRESS =  3'b010; 
localparam ADDRESS_ACK =    3'b011;
localparam WRITE_DATA =     3'b100;
localparam DATA_ACK =       3'b101;
localparam STOP =           3'b110;

reg         sda_out;
reg         scl_out;
reg [2:0]   counter = 0;
reg [7:0]   saved_addr;
reg [7:0]   saved_data;
reg         write;

reg [2:0]   current_state;
reg [2:0]   next_state;

assign sda_o = (write == 1) ? sda_out : 1;
assign scl_o = (write == 1) ? clk : 1;

// State register logic
always @(posedge clk, negedge rst_n) begin
    if (~rst_n)
        current_state <= IDLE;
    else
        current_state <= next_state;
end

// Counter logic
always @(posedge clk, negedge rst_n) begin
    if (current_state == WRITE_ADDRESS) begin
        counter <= counter - 1;
    end
    else if (current_state == WRITE_DATA) begin
        counter <= counter - 1;
    end 
end

// Next state combinational logic
always @* begin
    case (current_state)
        IDLE: begin
            if (enable) next_state = START;
            else        next_state = IDLE;
        end
        START:          next_state = WRITE_ADDRESS;
        WRITE_ADDRESS: begin
            if (counter == 0) begin
                        next_state = ADDRESS_ACK;
            end
        end
        ADDRESS_ACK:    next_state = WRITE_DATA;
        WRITE_DATA: begin
            if (counter == 0) begin
                        next_state = DATA_ACK;
            end
        end
        DATA_ACK:       next_state = STOP;
        default:        next_state = IDLE;
    endcase
end

// Output logic
always @(current_state, counter) begin
    case (current_state)
        IDLE: begin
            write       = 0;
            sda_out     = 1;
            scl_out     = 1;
            saved_addr  = {slave_address, rw};  // 1101.011.1
            saved_data  = {data_in};            // 1010.1010
        end
        START: begin
            sda_out     = 0;
            counter     = 7;
        end
        WRITE_ADDRESS: begin
            sda_out     = saved_addr[counter];
            write       = 1;
        end
        ADDRESS_ACK: begin
            write       = 0;
            sda_out     = 1;
            counter     = 7;
        end
        WRITE_DATA: begin
            write       = 1;
            sda_out     = saved_data[counter];
        end
        DATA_ACK: begin
            write       = 0;
            sda_out     = 1;
        end
        STOP: begin
            sda_out     = 1;
        end
    endcase
end
endmodule
