// Transmit slave address correctly
// Read 8 bytes from slave