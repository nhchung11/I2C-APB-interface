module TopLevel;
    reg clk 
endmodule