`ifndef SCOREBOARD
`define SCOREBOARD
   class scoreboard;
       bit [0:3] store;
   endclass
`endif